`timescale 1ps/1ps
module ROM (input [7:0] A,
            output [15:0] D);

    reg [15:0] rom [255:0];

    assign #10 D = rom[A];

    initial begin
        rom[0] = 16'b1001_110111111111;
        rom[1] = 16'b1001_001000001010;
        rom[2] = 16'b1010_111100000100;
        rom[3] = 16'b1010_000000000011;
        rom[4] = 16'b1001_010000000011;
        rom[5] = 16'b0110_010100100100;
        rom[6] = 16'b1100_000010010101;
        rom[7] = 16'b1001_000100000001;
        rom[8] = 16'b1110_000000001111;
        rom[9] = 16'b0100_110111010100;
        rom[10] = 16'b1111_001111111101;
        rom[11] = 16'b1111_001010001101;
        rom[12] = 16'b1111_000110011101;
        rom[13] = 16'b0000_100000100000;
        rom[14] = 16'b1001_011000000001;
        rom[15] = 16'b0100_001010000110;
        rom[16] = 16'b1010_111100000100;
        rom[17] = 16'b0000_100100010000;
        rom[18] = 16'b1001_010000000010;
        rom[19] = 16'b0100_001010000100;
        rom[20] = 16'b1010_111100000100;
        rom[21] = 16'b0000_000100011001;
        rom[22] = 16'b1000_111100111101;
        rom[23] = 16'b1000_100000101101;
        rom[24] = 16'b1000_100100011101;
        rom[25] = 16'b1001_010000000011;
        rom[26] = 16'b0000_110111010100;
        rom[27] = 16'b1110_000000001111;
    end

endmodule
